module test;


endmoule
